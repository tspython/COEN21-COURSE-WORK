module S0(A0,B0,F);
      input = A0, B0;
      output = F;
      assign F = A0 ^ B0;
end module